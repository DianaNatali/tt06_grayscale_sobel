`include "../src/parameters.svh" 

module sobel_control (
        input logic    clk_i,
        input logic    nreset_i,

        input logic    start_i,
        input logic    [PIXEL_WIDTH_OUT-1:0] in_px_gray_i,

        output logic   [PIXEL_WIDTH_OUT-1:0] out_px_sobel_o,
        output logic   px_ready_o
    );

    logic [SOBEL_COUNTER_MAX_BITS:0] counter_sobel;
    logic [MAX_RESOLUTION_BITS-1:0] counter_pixels;
    logic px_ready;
    
    sobel_matrix sobel_pixels; 

    logic [PIXEL_WIDTH_OUT-1:0] out_sobel_core;
    logic [PIXEL_WIDTH_OUT-1:0] out_sobel;

    typedef enum logic [2:0]{
        IDLE,
        FIRST_MATRIX, 
        NEXT_MATRIX, 
        END_FRAME} state_t;

    state_t fsm_state, next;

    sobel_core sobel(
        .matrix_pixels_i(sobel_pixels),
        .out_sobel_core_o(out_sobel_core)
    );


    always_ff @(posedge clk_i or negedge nreset_i)begin
        if(!nreset_i)begin
            fsm_state <= IDLE;
        end else begin
            fsm_state <= next;
        end
    end

    always_comb begin
        case(fsm_state)
            IDLE: begin
                if(start_i) next = FIRST_MATRIX;
                else next = IDLE;
            end
            FIRST_MATRIX: begin 
                if (counter_pixels == 1) next = NEXT_MATRIX; 
                else next = FIRST_MATRIX;
            end
            NEXT_MATRIX:begin
                if (start_i == 0) next = IDLE; 
                else next = NEXT_MATRIX;
            end
            default: next = IDLE;
        endcase
    end

    always_ff @(posedge clk_i or negedge nreset_i)begin
        if (!nreset_i)begin
            counter_sobel <= 'b0;
            counter_pixels <= 'b0;
            out_sobel <= 'b0;
            px_ready <= 'b0;
            sobel_pixels <= 'b0;
        end else begin
            case (next)
                IDLE: begin
                    px_ready <= 'b0;
                    out_sobel <= 'b0;
                    counter_pixels <= 'b0;
                    counter_sobel <= 'b0;
                end
                FIRST_MATRIX: begin
                    px_ready <= 'b0;
                    out_sobel <= '0;
                    case(counter_sobel)
                        1: sobel_pixels.vector0.pix0 <= in_px_gray_i;
                        2: sobel_pixels.vector0.pix1 <= in_px_gray_i;
                        3: sobel_pixels.vector0.pix2 <= in_px_gray_i;
                        4: sobel_pixels.vector1.pix0 <= in_px_gray_i;
                        5: sobel_pixels.vector1.pix1 <= in_px_gray_i;
                        6: sobel_pixels.vector1.pix2 <= in_px_gray_i;
                        7: sobel_pixels.vector2.pix0 <= in_px_gray_i;
                        8: sobel_pixels.vector2.pix1 <= in_px_gray_i;
                        9: sobel_pixels.vector2.pix2 <= in_px_gray_i;
                    endcase
                    counter_sobel <= counter_sobel + 1;
                    if (counter_sobel == 9) begin
                        counter_pixels <= counter_pixels + 1;
                        counter_sobel <= 'b0;
                        px_ready <= 'b1;
                        out_sobel <= out_sobel_core;
                        //out_sobel <= (out_sobel_core < SOBEL_THRESHOLD)? MIN_PIXEL_VAL : MAX_PIXEL_VAL-1;  //Binarization
                    end
                end
                NEXT_MATRIX: begin
                    px_ready <= 'b0;
                    out_sobel <= '0;
                    case(counter_sobel)
                        1: begin 
                            sobel_pixels.vector0 <= sobel_pixels.vector1;
                            sobel_pixels.vector1 <= sobel_pixels.vector2;
                            sobel_pixels.vector2.pix0 <= in_px_gray_i;
                        end
                        2: begin
                            sobel_pixels.vector2.pix1 <= in_px_gray_i;
                        end
                        3: begin
                            sobel_pixels.vector2.pix2 <= in_px_gray_i;
                        end
                    endcase
                    counter_sobel <= counter_sobel + 1;
                    if (counter_sobel == 3) begin
                        counter_pixels <= counter_pixels + 1;
                        counter_sobel <= 'b0;
                        px_ready <= 'b1;
                        out_sobel <= out_sobel_core;
                        //out_sobel <= (out_sobel_core < SOBEL_THRESHOLD)? MIN_PIXEL_VAL : MAX_PIXEL_VAL-1;  //Binarization
                    end
                end
                default: begin
                    px_ready <= 'b0;
                    out_sobel <= 'b0;
                    counter_pixels <= 'b0;
                    counter_sobel <= 'b0;
                end
            endcase
        end
    end


    assign  out_px_sobel_o = out_sobel;
    assign  px_ready_o = px_ready; 

endmodule
